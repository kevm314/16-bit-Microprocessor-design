LIBRARY ieee;
USE ieee.std_logic_1164.all;


ENTITY proc IS 
PORT (  
         SW : IN std_logic_vector(18 DOWNTO 0);
			LEDG: OUT std_logic_vector(15 DOWNTO 0);
			KEY: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			BusWires: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX3 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX4 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX5 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX6 : OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX7 : OUT STD_LOGIC_VECTOR(0 TO 6);
			Instructions : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			LEDR: OUT STD_LOGIC_VECTOR(16 DOWNTO 0));
END proc; 





ARCHITECTURE Behaviour OF proc IS


--register final hex outputs

SIGNAL hexin: STD_LOGIC_VECTOR(15 downto 0);
SIGNAL hexin2: STD_LOGIC_VECTOR(15 downto 0);

SIGNAL dummy: STD_LOGIC_VECTOR(15 DOWNTO 0);

--ALUdata output
SIGNAL ALUdata1 : STD_LOGIC_VECTOR(15 DOWNTO 0); 
SIGNAL Karry : STD_LOGIC ;



-- main input into the Control Unit via the processorSIGNAL Reset : STD_LOGIC;
SIGNAL wCu : STD_LOGIC;SIGNAL CLoK : STD_LOGIC;SIGNAL F : STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL PDone : STD_LOGIC;

  --  driving signals for register entering and exiting data
SIGNAL RProin, RProout : STD_LOGIC_VECTOR(7 DOWNTO 0); 

TYPE Rdata IS ARRAY (7 downto 0) OF std_logic_vector(15 downto 0);
SIGNAL RDAT : Rdata;

  -- to enable data to enter register
SIGNAL APin, GPin, GPout : STD_LOGIC;

 -- actual register data that will exit
SIGNAL Adata, Gdata, Idata, instruction : STD_LOGIC_VECTOR(15 DOWNTO 0);

-- actual external data signals
SIGNAL Data : STD_LOGIC_VECTOR(15 DOWNTO 0);


-- control signals for external data and ALU
SIGNAL Extern : STD_LOGIC ;
SIGNAL AddSub : STD_LOGIC_VECTOR(1 DOWNTO 0); -- function and register operand signals from instruction registerSIGNAL F: STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL REX, REY : STD_LOGIC_VECTOR(2 DOWNTO 0); 
-- program address as generated by the program counter
SIGNAL PROGcount : std_logic_vector(7 downto 0);

SIGNAL isInstruction : STD_LOGIC;

--RAM
COMPONENT progMem16 IS
GENERIC ( S : INTEGER := 16;
	N : INTEGER := 8 );
port(
	clock : in std_logic; -- brought in from the processor
	data_in : in std_logic_vector (15 downto 0); -- this is not required
	write_addr : in std_logic_vector (N-1 downto 0); -- this is not required
	read_addr : in std_logic_vector (N-1 downto 0); -- this is brought in from the program counter
	write_enable : in std_logic; --this always 1
	data_out : out std_logic_vector (15 downto 0)); --this links to external in
END COMPONENT;





--the program counter
COMPONENT programCounter IS 
PORT (	       
					cluk : IN std_logic; --clock
				 specify: IN std_logic_vector(7 downto 0); --specific address to count from
		 resetCounter : IN std_logic; -- to reset must pass 00000000 as the specify address
		  enableCount : IN std_logic; --variable to enable counting
				  count : OUT std_logic_vector(7 downto 0)); --the actual output address to be used by RAM
END COMPONENT; 







 -- n-bit adder/sub
COMPONENT myALU IS 
PORT (	        A : IN std_logic_vector(15 downto 0);
                 B : IN std_logic_vector(15 downto 0); 
                 As: IN std_logic_vector(1 downto 0); --As is AddSub signal control signal
                 G : OUT std_logic_vector(15 downto 0);
	          Kcarry: OUT std_logic);
END COMPONENT;


 --control unit
COMPONENT controlunit IS
PORT (	       
	     w : IN std_LOGIC;
	  clock: IN std_logic;
       Fcu: IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- 3 instruction bits
		 Rx : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Rx 3 bits from instruction
		 Ry : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Ry 3 bits from instruction
		 Rin: OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --driving ENTERING data for all registers
		Rout: OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --driving EXITING data for all registers VIA A MULTIPLEXER OR TRINODE STRUCTURE
       Ain: OUT std_logic;
	    Gin: OUT std_logic;
	   Gout: OUT std_logic;
 AddSubXOR: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
  ExternIn: OUT std_logic;
		 isI: OUT std_logic;
	   Done: OUT std_logic);
END COMPONENT;



--16 bit register
--component structure for proc hierarchy
COMPONENT R16bReg IS 
	PORT (
       Dreg : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	       clk : IN STD_LOGIC;
      enable: IN STD_LOGIC;
	      Qreg: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));        
END COMPONENT;


--trinode buffer
COMPONENT tristate is
  port( 		    Atr : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				 enable : in std_logic;
                Qtr : out std_logic_VECTOR(15 DOWNTO 0));
end COMPONENT;


--hexdecode
COMPONENT hexdecode is
	port ( A : IN std_logic_vector(3 downto 0);
			D : OUT std_logic_vector(0 to 6));
end COMPONENT;

BEGIN


-- redirect inputs to control signals
CLoK <= KEY(0);
wCu <= SW(17);
--HEX0(0 TO 6) <= PROGcount(6 DOWNTO 0);
--instruction <= SW(15 DOWNTO 0);
instruction <= DATA;

Instructions <= instruction;

F <= Idata(15 DOWNTO 13);
REX <= Idata(12 DOWNTO 10);
REY <= Idata(9 DOWNTO 7);

--redirect control signals to outputs
--LEDR(15 DOWNTO 0) <= BusWires;




-- generate code for 8 general purpose registers and A, G registers

-- 8 GPR
-- signals to be defined BusWires, RegIn(15 to 0), RegOut(15 to 0)

gpr: FOR i IN 7 DOWNTO 0 GENERATE

	FA0: R16bReg port map(BusWires, CLoK, RProin(i), RDAT(i));
	MainRegisters: tristate port map(RDAT(i), RProout(i), BusWires);

END GENERATE gpr;
--export data through trinode structure



--A and G and instruction registers

Areg: R16bReg port map(BusWires, CLoK, APin, Adata);

-- Gdata output driven to bus via a trinode buffer using GPout
Greg: R16bReg port map(ALUdata1, CLoK, GPin, Gdata); 
Gregister: tristate port map(Gdata, GPout, BusWires);


--data external input
Externally: tristate port map(Data, Extern, BusWires);





-- Instruction register
Ireg: R16bReg port map(instruction, CLoK, isInstruction, Idata); 


-- Mapping to control unit through instruction register signals and other control signals

CU: controlunit port map (wCu, CLoK, F, REX, REY, RProin, RProout, APin, GPin, GPout, AddSub, Extern, isInstruction, PDone);
AluSection: myALU port map (Adata, BusWires, AddSub, ALUdata1, Karry);



--hexin <= RDAT(1) WHEN KEY(1)='0' ELSE
--RDAT(2) WHEN KEY(2)='0' ELSE
--RDAT(3) WHEN KEY(3)='0' ELSE RDAT(0);


--hexin2 <= RDAT(5) WHEN KEY(1)='0' ELSE
--RDAT(6) WHEN KEY(2)='0' ELSE
--RDAT(7) WHEN KEY(3)='0' ELSE RDAT(4);

--test the first two registers
hexin <= RDAT(0);
hexin2 <= RDAT(1);

h3: hexdecode port map (hexin(15 downto 12), hex3);
h2: hexdecode port map (hexin(11 downto 8), hex2);
h1: hexdecode port map (hexin(7 downto 4), hex1);
h0: hexdecode port map (hexin(3 downto 0), HEX0);


h7: hexdecode port map (hexin2(15 downto 12), hex7);
h6: hexdecode port map (hexin2(11 downto 8), hex6);
h5: hexdecode port map (hexin2(7 DOWNTO 4), hex5);
h4: hexdecode port map (hexin2(3 downto 0), hex4);


--RAM and program Counter

vRam: progMem16 port map (CLoK, "0000000000000111", "00000000", PROGcount, '0', DATA);
ProgC: programCounter port map (PDone, "00000000", NOT wCu, '1', PROGcount); --2nd last is enable count, 3rd last is official reset

dummy <= RDAT(0);

LEDG(15 DOWNTO 0) <= RDAT(0)(15 DOWNTO 0);
LEDR(15 DOWNTO 0) <= BusWires;
LEDR(16) <= PDone;				  
				  
				  
END Behaviour;

